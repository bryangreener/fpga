module top(
	input logic clk, //100MHz
	output logic led
);
endmodule