module fp_add (
    input clk,
    input rst,
    input [31:0] a,
    input [31:0] b,
    output [31:0] c
);


endmodule